

/*
	Bit 5 in the SREG in NOT implemented (Half carry)

*/

module BasicMCUInFPGA(input clk,
							output [15:0]digitalIO,
							output stuck,
							input butt,
							output [7:0]debug,
							input RXD,
							input buttProg,
							input reset,
							output progMode);

assign stuck=(state==STUCK);

assign progMode=programmingMode;

assign digitalIO=(programmingMode==1'b1)?8'b10101010:{3'd0,IOregs[8'd5][5:0],IOregs[8'd11]};

//assign digitalIO={flash_out_1,flash_out_2};
//assign digitalIO=(buttProg==1'b1)?{flash_out_1}:nextByteProgCounter;
//assign digitalIO={8'd0,OPCODE};	
//assign digitalIO=readdata;
//assign digitalIO={IOregs[62],reg1output};
assign debug={OPCODE[3:0],state};	
				
				
//Register file
reg [7:0]reg1input;
reg writeEn;
reg [4:0]reg1address;
wire [7:0]reg1output;

reg [7:0]reg2address;
wire [7:0]reg2output;

reg [7:0]SREG;

reg [15:0]SP;
reg [13:0]RA;

reg [15:0]PC;

reg [7:0]IOregs[64];


//Flash
reg [13:0]flash_addr_1;
reg [13:0]flash_addr_2;

reg [15:0]flash_dataIN_1;
reg [15:0]flash_dataIN_2;
reg flash_WRen_1;
wire flash_WRen_2;

assign flash_WRen_2=0;

wire [15:0]flash_out_1;
wire [15:0]flash_out_2;

//RAM
reg [10:0]ram_address;
reg [7:0]ram_inputData;
wire [7:0]ram_outputData;
reg ram_WRen;


//Working regs
reg [3:0]state;
parameter FETCH=4'd0,FETCH2=4'd1,FETCH3=4'd2,WORK1=4'd3,WORK2=4'd4,WORK3=4'd5,STUCK=4'd6;

reg [15:0]readedByte1;
reg [15:0]readedByte2;

wire [7:0]OPCODE;

localparam error=8'd0,
ldi=8'd1,
jmp=8'd2,
call=8'd3,
out=8'd4,
ret=8'd5,
cli=8'd6,
rjmp=8'd7,
eor=8'd8,
subi=8'd9,
sbci=8'd10,
brne=8'd11,
nop=8'd12;	

wire finalClock;
wire slowclk;

assign finalClock=clk;

slowClock cloco(clk, slowclk);



wire [7:0]readdata;
wire dataCount;
UART prog(readdata,dataCount,RXD,clk);


instructionSelector selector(readedByte1,OPCODE);


wire myClock;

PushButton_Debouncer debouncer(slowClock,butt,myClock);


registerFile regFile(finalClock,reg1input,writeEn,reg1address,reg1output,reg2address,reg2output);

FLASH flash((programmingMode==1'b0)?PC:flash_addr_1,PC+1,finalClock,flash_dataIN_1,flash_dataIN_2,flash_WRen_1,flash_WRen_2,flash_out_1,flash_out_2);
//FLASH flash(PC,PC+1,finalClock,flash_dataIN_1,flash_dataIN_2,flash_WRen_1,flash_WRen_2,flash_out_1,flash_out_2);


RAM ram(ram_address,finalClock,ram_inputData,ram_WRen,ram_outputData);

reg programmingMode;



always @(posedge finalClock)
begin
		
	if(programmingMode==1'b0)
	begin
		case (state)
				
		FETCH:
		begin
			//Wait for the RAM to output the data			
			state=FETCH2;
		end
		
		FETCH2:
		begin
			readedByte1={flash_out_1[7:0],flash_out_1[15:8]}; //Read PC
			readedByte2={flash_out_2[7:0],flash_out_2[15:8]}; //Read PC+1 (For 32bit instructions
			//state=WORK1; //Set the state to work
		//	PC=PC+1;
			state=FETCH3;
		end
		
		FETCH3:
		begin //The instructionSelector does its job in this tick
			state=WORK1;
		end
		
		WORK1:
		begin
			
			case (OPCODE)
				ldi: 
				begin
					reg1address=5'd16+readedByte1[7:4]; //Calculates the register to write the info to
					reg1input={readedByte1[11:8],readedByte1[3:0]};
					writeEn=1'b1; 
					//Go to next state now,while the value is being stored
				end
				
				
				jmp:
				begin
					PC={readedByte2[15:0]}; //Set new value for PC (We are not using the full 32 bit as the datasheet seys (we don't need it for the ATMega328P
				end
				
				
				call:
				begin
					//Store to the stack the next address										
					ram_address=SP; //Store the next instruction into the address
					PC=PC+16'd2; //Sets the PC to the next instruction, to save to the stack this value
					ram_inputData=PC[15:8]; //Save the most significant digits to the first stack
					ram_WRen=1'b1;
					//Go to the next state by default, while the data1 is stored
				end
				
				
				out:
				begin
					writeEn=1'b0; //Just in case, we sent writeEn to 0
					reg1address=readedByte1[8:4]; //Request the data in the register file stored in the register we want
					//Wait just in case the register file taskes 1 cycle to output the data
				end
				
				ret:
				begin
					SP=SP+14'd2; //Increment the stack by 2
					ram_WRen=1'b0; //Make sure we are not writing
					ram_address=SP; //Set the stack address to read
					//Waits for the ram to provide the data
					state=WORK2;
				end
			
				
				cli:
				begin
					SREG[7]=1'b0;  //Disable interrupt pin
					PC=PC+16'd1;
				end
			
				rjmp:
				begin
					PC=PC+({readedByte1[11],readedByte1[11],readedByte1[11],readedByte1[11],readedByte1[11:0]})+16'd1;  //Jump to the sign extended offset +1
				end
				
				eor:
				begin				
					writeEn=1'b0;  //Make sure we are not writing					
					reg1address=readedByte2[8:4]; //Read r1
					reg2address={readedByte1[9],readedByte1[3:0]}; //Read r2
					//Wait just in case for the register file
				end
				
				
				subi:
				begin
					writeEn=1'b0; //We are reading 
					reg1address=5'd16+readedByte1[7:4];  //Register we are substracing from and to (16-32)
					//Wait until next cycle for the output
				end
				
				sbci:
				begin
					writeEn=1'b0; //We are reading 
					reg1address=5'd16+readedByte1[7:4];  //Register we are substracing from and to (16-32)
					//Wait until next cycle for the output
				end
				
				brne:
				begin
					if(SREG[1]==1'b0) //If the zero flag is NOT set (Not equal), branch
					begin
						PC=PC+({readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9],readedByte1[9:3]})+16'd1;  //Jump to the sign extended offset +1				
					end
					else
					begin
						PC=PC+16'd1;
					end				
				end
				
				nop:
				begin
					
				end	
				
			endcase
	
			if(OPCODE==error) state=STUCK;
			else state=WORK2;
			
		end
		
		WORK2:
		begin
		
			case (OPCODE)
				ldi: 
				begin					
					//The value should be stored now,finish the instruction
					writeEn=1'b0; //Disable the writeEnable for the register file
					PC=PC+16'd1;					
				end	
				
				call:
				begin
					//Store to the stack the next address										
					ram_address=SP-14'b1; //Store the next instruction into the address				
					ram_inputData=PC[7:0]; //Save the LEAST significant digits to the first stack
					ram_WRen=1'b1;
					//Go to the next state by default, while the data2 is stored				
				end
				
				
				out:
				begin
					IOregs[{readedByte1[10:9],readedByte1[3:0]}]=reg1output;  //Set the right IO register to the data in the register file output
					if({readedByte1[10:9],readedByte1[3:0]}==6'b111101) SP[7:0]=reg1output;  //If the IO reg is 61, it is SPl
					if({readedByte1[10:9],readedByte1[3:0]}==6'b111110) SP[15:8]=reg1output; //If the IO reg is 62, its is SPH
					PC=PC+16'd1;		
				end
				
				ret:
				begin
					PC[7:0]=ram_outputData; //Set the MSB of the PC to the data from the stack
					ram_address=SP-14'b1; //Read the LSB part
					//Wait until the LSB part can be read
				end	
				
				eor:
				begin
				   reg1input=reg1output^reg2output; //Do the xor operation and store it in the first register					
					writeEn=1'b1; //Enable the writing
					//Wait for the write
				end
							
			
				subi:
				begin
					//Address should already be set from the last step
					reg1input=reg1output-{readedByte1[11:8],readedByte1[3:0]};
					SREG[3]=(reg1output[7] & !readedByte1[11] & !reg1input[7])|(!reg1output[7] & readedByte1[11] & reg1input[7]);
					SREG[0]= (!reg1output[7] & readedByte1[11])|(readedByte1[11] & reg1input[7])|(reg1input[7] & !reg1output[7]);	
					writeEn=1'b1; 
					//Go to next state now,while the value is being stored
				end
				
				sbci:
				begin
					//Address should already be set from the last step
					reg1input=reg1output-{readedByte1[11:8],readedByte1[3:0]}-SREG[0];
					SREG[3]=(reg1output[7] & !readedByte1[11] & !reg1input[7])|(!reg1output[7] & readedByte1[11] & reg1input[7]);
					SREG[0]= (!reg1output[7] & readedByte1[11])|(readedByte1[11] & reg1input[7])|(reg1input[7] & !reg1output[7]);	
					writeEn=1'b1; 
					//Go to next state now,while the value is being stored
				end				
				
			endcase			
			
			state=WORK3;
		end
		
		WORK3:
		begin
			case (OPCODE)
			
				call:
				begin		
					ram_WRen=1'd0;  //Stop writing to the ram
					PC={readedByte1[8:4],readedByte1[0],readedByte2[15:0]};  //Go to the address in the instruction					
					SP=SP-14'd2; //Decrease the stack pointer by 2 (Its is a postdecrement)
					//Finished, go on with the execution					
				end
					
				ret:
				begin
					PC[15:8]=ram_outputData; //Set the MSB of the PC to the data from the stack
					//Finished, go on with the execution				
				end
				
				eor:
				begin
					writeEn=1'b0; //Disable writing to the register file
					SREG[3]=1'b0;
					SREG[2]=reg1input[7];					
					SREG[1]=(reg1input==8'b0);					
					PC=PC+16'd1;
					//Finished, go on with the execution	
				end	
			
				subi:
				begin					
					writeEn=1'b0;  //Disable writing	
					SREG[2]=reg1input[7];					
					SREG[1]=(reg1input==8'b0);	
					PC=PC+16'd1;
					//Finished, go on with the execution				
				end
				
				sbci:
				begin					
					writeEn=1'b0;  //Disable writing	
					SREG[2]=reg1input[7];					
					SREG[1]=(reg1input==8'b0) & SREG[1];	 //Keeps the old value unless the result is not 0
					PC=PC+16'd1;
					//Finished, go on with the execution				
				end
				
				nop:
				begin
					PC=PC+16'd1;					
				end
					
			
			endcase			
			
			state=FETCH;
		end
		
		STUCK:
		begin
			//Stay here until the Wraiths destroy this planet :P
		end
		
	endcase
	
	SREG[4]=SREG[3]^SREG[2]; //Update the XOR in the SREG register
	
	IOregs[61]=SP[7:0];   //Update real IO stack registers from the SP that we use
	IOregs[62]=SP[15:8];
	
	flash_WRen_1=0;
	case(progDetect)
	4'd0:
	begin
		if(readdata==8'd169) progDetect=4'd1;
	end
	4'd1:
	begin
		if(readdata==8'd68) progDetect=4'd2;
	end
	4'd2:
	begin
		if(readdata==8'd69) 
		begin
			programmingMode=1'b1;
			lastRXstate=dataCount;
			nextByteProgCounter=0;
			timeToExitProgramming=40'd5000000;
			progDetect=4'd0;			
		end
	end
	default:
	begin
		progDetect=4'd0;
	end
	endcase
	
	
	end
	else 
	begin
			
		if(lastRXstate!=dataCount)
		begin
			timeToExitProgramming=40'd5000000;
			if(nextByteProgCounter%2==0)
			begin
				flash_WRen_1=0;
				flash_dataIN_1[15:8]=readdata;
				flash_addr_1=nextByteProgCounter/2;
			end
			else
			begin
				flash_WRen_1=1;
				flash_dataIN_1[7:0]=readdata;

			end				
			
			nextByteProgCounter=nextByteProgCounter+1;
			lastRXstate=dataCount;							
		end
		else 
		begin
			timeToExitProgramming=timeToExitProgramming-1;
			if(timeToExitProgramming<=0)
			begin
				 programmingMode=0;
				flash_WRen_1=0;
			end
		end
		
		
		PC=0;
		SP=0;
		SREG=0;
		state=FETCH;
		IOregs[8'd5]=0;
		IOregs[8'd11]=0;
	end
	
end


reg [49:0]nextByteProgCounter;
reg lastRXstate;

reg [3:0]progDetect;


reg [39:0]timeToExitProgramming;




endmodule